efwef
sdfwef

  jhgdsfjwsekfhwe
