efwef
sdfwef
